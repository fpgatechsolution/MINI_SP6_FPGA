
----------------------------------------------------------------------------------
-- COMPANY      : FPGATECHSOLUTION
-- MODULE NAME  : UART_RECEIVER
-- URL     		: WWW.FPGATECHSOLUTION.COM
----------------------------------------------------------------------------------
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY TOP IS
    PORT ( 
		CLOCK_12MHZ : IN  STD_LOGIC;
		
    	LED_RED  	: OUT  STD_LOGIC;
		LED_GREEN 	: OUT  STD_LOGIC;
		LED_BLUE 	: OUT  STD_LOGIC;
		
		PUSH_BTN_1 	: IN  STD_LOGIC;
		PUSH_BTN_2 	: IN  STD_LOGIC;
		PUSH_BTN_3 	: IN  STD_LOGIC;
		PUSH_BTN_4 	: IN  STD_LOGIC;

		DIP_SW_1	: IN  STD_LOGIC;
		DIP_SW_2	: IN  STD_LOGIC;
		DIP_SW_3	: IN  STD_LOGIC;
		DIP_SW_4	: IN  STD_LOGIC;
		
		LED			: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        
		USB_UART_RX : IN  STD_LOGIC;
        USB_UART_TX : OUT  STD_LOGIC;
		
		IO_J1_3  	: OUT STD_LOGIC;
		IO_J1_4  	: OUT STD_LOGIC;
		IO_J1_5  	: OUT STD_LOGIC;
		IO_J1_6  	: OUT STD_LOGIC;
		IO_J1_7  	: OUT STD_LOGIC;
		IO_J1_8  	: OUT STD_LOGIC;
		IO_J1_9  	: OUT STD_LOGIC;
		IO_J1_10  	: OUT STD_LOGIC;
		IO_J1_11	: OUT STD_LOGIC;
		IO_J1_12	: OUT STD_LOGIC;
		IO_J1_13	: OUT STD_LOGIC;
		IO_J1_14	: OUT STD_LOGIC;
		IO_J1_15	: OUT STD_LOGIC;
		IO_J1_16	: OUT STD_LOGIC;
		IO_J1_17	: OUT STD_LOGIC;
		IO_J1_18	: OUT STD_LOGIC;
		IO_J1_19	: OUT STD_LOGIC;
		IO_J1_20	: OUT STD_LOGIC;
		IO_J1_21	: OUT STD_LOGIC;
		IO_J1_22	: OUT STD_LOGIC;
		IO_J1_23	: OUT STD_LOGIC;
		IO_J1_24	: OUT STD_LOGIC;
		IO_J1_25	: OUT STD_LOGIC;
		IO_J1_26	: OUT STD_LOGIC;
		IO_J1_27	: OUT STD_LOGIC;
		IO_J1_28	: OUT STD_LOGIC;
		IO_J1_29	: OUT STD_LOGIC;
		IO_J1_30	: OUT STD_LOGIC;
		IO_J1_31	: OUT STD_LOGIC; 
		IO_J1_32	: OUT STD_LOGIC;
		IO_J1_33	: OUT STD_LOGIC;
		IO_J1_35	: OUT STD_LOGIC;
		IO_J1_36	: OUT STD_LOGIC;
		IO_J1_37	: OUT STD_LOGIC;
		IO_J1_38	: OUT STD_LOGIC;
	
		IO_J2_3 	: OUT STD_LOGIC;
		IO_J2_4 	: OUT STD_LOGIC;
		IO_J2_5 	: OUT STD_LOGIC;
		IO_J2_6 	: OUT STD_LOGIC;
		IO_J2_7 	: OUT STD_LOGIC;
		IO_J2_8 	: OUT STD_LOGIC;
		IO_J2_9 	: OUT STD_LOGIC;
		IO_J2_10	: OUT STD_LOGIC;
		IO_J2_11	: OUT STD_LOGIC;
		IO_J2_12	: OUT STD_LOGIC;
		IO_J2_13	: OUT STD_LOGIC;
		IO_J2_14	: OUT STD_LOGIC;
		IO_J2_15	: OUT STD_LOGIC;
		IO_J2_16	: OUT STD_LOGIC;
		IO_J2_17	: OUT STD_LOGIC;
		IO_J2_18	: OUT STD_LOGIC;
		IO_J2_19	: OUT STD_LOGIC;
		IO_J2_20	: OUT STD_LOGIC;
		IO_J2_21	: OUT STD_LOGIC;
		IO_J2_22	: OUT STD_LOGIC;
		IO_J2_23	: OUT STD_LOGIC;
		IO_J2_24	: OUT STD_LOGIC;
		IO_J2_25	: OUT STD_LOGIC;
		IO_J2_26	: OUT STD_LOGIC;
		IO_J2_27	: OUT STD_LOGIC;
		IO_J2_28	: OUT STD_LOGIC;
		IO_J2_29	: OUT STD_LOGIC;
		IO_J2_30	: OUT STD_LOGIC;
		IO_J2_31	: OUT STD_LOGIC;
		IO_J2_32	: OUT STD_LOGIC;
		IO_J2_33	: OUT STD_LOGIC;
		IO_J2_34	: OUT STD_LOGIC;
		IO_J2_35	: OUT STD_LOGIC;
		IO_J2_36	: OUT STD_LOGIC;
		IO_J2_37	: OUT STD_LOGIC;
		IO_J2_38	: OUT STD_LOGIC

);
END TOP;

ARCHITECTURE BEHAVIORAL OF TOP IS

	COMPONENT UART_CONTROL
		PORT(
			RESET : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			RXD : IN STD_LOGIC;          
			TXD : OUT STD_LOGIC;
			TEST_LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
			);
	END COMPONENT;


	COMPONENT LED_SHIFTER
		PORT(
			SEL : IN STD_LOGIC;   
			INDX : IN STD_LOGIC_VECTOR(3 DOWNTO 0);          
			LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
			);
	END COMPONENT;

SIGNAL COUNT_RGB : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LED_RX    : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LED_SHIFT : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COUNT   	 : STD_LOGIC_VECTOR(23 DOWNTO 0); 
SIGNAL CLK_1S	 : STD_LOGIC;

BEGIN

	INST_UART_CONTROL: UART_CONTROL PORT MAP(
		RESET 	=>PUSH_BTN_2 ,
		CLK   	=>CLOCK_12MHZ ,
		RXD   	=>USB_UART_RX ,
		TXD      =>USB_UART_TX ,
		TEST_LED=> LED_RX
	);




	PROCESS (CLOCK_12MHZ) 
		BEGIN
			IF PUSH_BTN_1='1'  THEN 
				COUNT <= (OTHERS => '0');
			ELSIF CLOCK_12MHZ='1' AND CLOCK_12MHZ'EVENT THEN
				COUNT <= COUNT + 1;
			END IF;
	END PROCESS;
	
	CLK_1S<=COUNT(22);
	
	PROCESS (CLK_1S) 
		BEGIN
			IF PUSH_BTN_1='1'  THEN 
				COUNT_RGB <= (OTHERS => '0');
			ELSIF CLK_1S='1' AND CLK_1S'EVENT THEN
				COUNT_RGB <= COUNT_RGB + 1;
			END IF;
	END PROCESS;
	


	  
    LED_RED <=COUNT_RGB(0) WHEN (DIP_SW_1='0') ELSE (PUSH_BTN_1 OR PUSH_BTN_2 OR PUSH_BTN_3 OR PUSH_BTN_4) ;
    LED_GREEN<=COUNT_RGB(1) WHEN (DIP_SW_1='0') ELSE (DIP_SW_2 OR DIP_SW_3 OR DIP_SW_4 ) ;
    LED_BLUE<=COUNT_RGB(2); 

LED<=LED_SHIFT WHEN (DIP_SW_1='0') ELSE LED_RX;

	INST_LED_SHIFTER: LED_SHIFTER 
	PORT MAP
		(
			SEL=>DIP_SW_4,
			INDX =>COUNT_RGB(3 DOWNTO 0) ,
			LED => LED_SHIFT
		);


	LED<=LED_SHIFT WHEN (DIP_SW_1='0') ELSE LED_RX;
	
	
	IO_J1_3	 <=DIP_SW_3;
	IO_J1_4	 <=DIP_SW_3; 
	IO_J1_5	 <=DIP_SW_3; 
	IO_J1_6	 <=DIP_SW_3; 
	IO_J1_7	 <=DIP_SW_3; 
	IO_J1_8	 <=DIP_SW_3; 
	IO_J1_9  <=DIP_SW_3; 
	IO_J1_10 <=DIP_SW_3; 
	IO_J1_11 <=DIP_SW_3; 
	IO_J1_12 <=DIP_SW_3; 
	IO_J1_13 <=DIP_SW_3; 
	IO_J1_14 <=DIP_SW_3; 
	IO_J1_15 <=DIP_SW_3; 
	IO_J1_16 <=DIP_SW_3; 
	IO_J1_17 <=DIP_SW_3; 
	IO_J1_18 <=DIP_SW_3; 
	IO_J1_19 <=DIP_SW_3; 
	IO_J1_20 <=DIP_SW_3; 
	IO_J1_21 <=DIP_SW_3; 
	IO_J1_22 <=DIP_SW_3; 
	IO_J1_23 <=DIP_SW_3; 
	IO_J1_24 <=DIP_SW_3; 
	IO_J1_25 <=DIP_SW_3; 
	IO_J1_26 <=DIP_SW_3; 
	IO_J1_27 <=DIP_SW_3; 
	IO_J1_28 <=DIP_SW_3; 
	IO_J1_29 <=DIP_SW_3; 
	IO_J1_30 <=DIP_SW_3; 
	IO_J1_31 <=DIP_SW_3; 
	IO_J1_32 <=DIP_SW_3; 
	IO_J1_33 <=DIP_SW_3; 
	IO_J1_35 <=DIP_SW_3; 
	IO_J1_36 <=DIP_SW_3; 
	IO_J1_37 <=DIP_SW_3; 
	IO_J1_38 <=DIP_SW_3; 
	
	IO_J2_3  <=DIP_SW_3; 
	IO_J2_4  <=DIP_SW_3; 
	IO_J2_5  <=DIP_SW_3; 
	IO_J2_6  <=DIP_SW_3; 
	IO_J2_7  <=DIP_SW_3; 
	IO_J2_8  <=DIP_SW_3; 
	IO_J2_9  <=DIP_SW_3; 
	IO_J2_10 <=DIP_SW_3; 
	IO_J2_11 <=DIP_SW_3; 
	IO_J2_12 <=DIP_SW_3; 
	IO_J2_13 <=DIP_SW_3; 
	IO_J2_14 <=DIP_SW_3; 
	IO_J2_15 <=DIP_SW_3; 
	IO_J2_16 <=DIP_SW_3; 
	IO_J2_17 <=DIP_SW_3; 
	IO_J2_18 <=DIP_SW_3; 
	IO_J2_19 <=DIP_SW_3; 
	IO_J2_20 <=DIP_SW_3; 
	IO_J2_21 <=DIP_SW_3; 
	IO_J2_22 <=DIP_SW_3; 
	IO_J2_23 <=DIP_SW_3; 
	IO_J2_24 <=DIP_SW_3; 
	IO_J2_25 <=DIP_SW_3; 
	IO_J2_26 <=DIP_SW_3; 
	IO_J2_27 <=DIP_SW_3; 
	IO_J2_28 <=DIP_SW_3; 
	IO_J2_29 <=DIP_SW_3; 
	IO_J2_30 <=DIP_SW_3; 
	IO_J2_31 <=DIP_SW_3; 
	IO_J2_32 <=DIP_SW_3; 
	IO_J2_33 <=DIP_SW_3; 
	IO_J2_34 <=DIP_SW_3; 
	IO_J2_35 <=DIP_SW_3; 
	IO_J2_36 <=DIP_SW_3; 
	IO_J2_37 <=DIP_SW_3; 
	IO_J2_38 <=DIP_SW_3; 
	
	

END BEHAVIORAL;

