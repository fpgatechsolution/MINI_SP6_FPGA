
----------------------------------------------------------------------------------
-- COMPANY      : FPGATECHSOLUTION
-- MODULE NAME  : UART_RECEIVER
-- URL     		: WWW.FPGATECHSOLUTION.COM
----------------------------------------------------------------------------------
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY TOP IS
    PORT ( 
		CLOCK_100MHZ : IN  STD_LOGIC;
        RESET_n: IN  STD_LOGIC;
		
		RGB_LED1: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		RGB_LED2: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        
		USB_UART_RX : IN  STD_LOGIC;
        USB_UART_TX : OUT  STD_LOGIC
		


);
END TOP;

ARCHITECTURE BEHAVIORAL OF TOP IS

	COMPONENT UART_CONTROL
		PORT(
			RESET : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			RXD : IN STD_LOGIC;          
			TXD : OUT STD_LOGIC;
			TEST_LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
			);
	END COMPONENT;


	COMPONENT LED_SHIFTER
		PORT(
			SEL : IN STD_LOGIC;   
			INDX : IN STD_LOGIC_VECTOR(3 DOWNTO 0);          
			LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
			);
	END COMPONENT;


	COMPONENT dcm_wrapper
		PORT(
			sys_clock : IN STD_LOGIC;          
			clk_out12 : OUT STD_LOGIC
			);
	END COMPONENT;
	
	
SIGNAL COUNT_RGB : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LED_RX    : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LED_SHIFT : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COUNT   	 : STD_LOGIC_VECTOR(23 DOWNTO 0); 
SIGNAL CLK_1S	 : STD_LOGIC;

SIGNAL CLOCK_12MHZ: STD_LOGIC;
SIGNAL RESET: STD_LOGIC;

BEGIN


RESET<= NOT RESET_n;

INST_dcm_wrapper: dcm_wrapper PORT MAP(
		sys_clock 	=>CLOCK_100MHZ ,
		clk_out12   =>CLOCK_12MHZ);



	INST_UART_CONTROL: UART_CONTROL PORT MAP(
		RESET 	=> RESET ,
		CLK   	=>CLOCK_12MHZ ,
		RXD   	=>USB_UART_RX ,
		TXD      =>USB_UART_TX ,
		TEST_LED=> LED_RX
	);




	PROCESS (CLOCK_12MHZ) 
		BEGIN
			IF RESET='1'  THEN 
				COUNT <= (OTHERS => '0');
			ELSIF CLOCK_12MHZ='1' AND CLOCK_12MHZ'EVENT THEN
				COUNT <= COUNT + 1;
			END IF;
	END PROCESS;
	
	CLK_1S<=COUNT(22);
	
	PROCESS (CLK_1S) 
		BEGIN
			IF RESET='1'  THEN 
				COUNT_RGB <= (OTHERS => '0');
			ELSIF CLK_1S='1' AND CLK_1S'EVENT THEN
				COUNT_RGB <= COUNT_RGB + 1;
			END IF;
	END PROCESS;
	


	  



	INST_LED_SHIFTER: LED_SHIFTER 
	PORT MAP
		(
			SEL=>'1',
			INDX =>COUNT_RGB(3 DOWNTO 0) ,
			LED => LED_SHIFT
		);


	RGB_LED1<=NOT (LED_SHIFT(2 DOWNTO 0));
	RGB_LED2<=NOT (LED_SHIFT(5 DOWNTO 3)) ;
	

	
	

END BEHAVIORAL;

