----------------------------------------------------------------------------------
-- COMPANY      : FPGATECHSOLUTION
-- MODULE NAME  : UART_TRANSMITTER
-- URL     		: WWW.FPGATECHSOLUTION.COM
----------------------------------------------------------------------------------
--


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY UART_TRANSMITTER IS
	GENERIC
	(
		FREQUENCY	: INTEGER;
		BAUD		: INTEGER
	);
	PORT
	(
		CLK			: IN STD_LOGIC;
		TXD			: OUT STD_LOGIC;
		TXD_DATA	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		TXD_START	: IN STD_LOGIC;
		TXD_BUSY	: OUT STD_LOGIC
	);
END ENTITY UART_TRANSMITTER;

ARCHITECTURE TRANSMITTER_BEH OF UART_TRANSMITTER IS

TYPE STATE_TYPE IS (IDLE, START, BIT0, BIT1, BIT2, BIT3, BIT4, BIT5, BIT6, BIT7, STOP1, STOP2);

SIGNAL STATE : STATE_TYPE := IDLE; 
SIGNAL DATA : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL BAUD_TICK : STD_LOGIC;
SIGNAL BUSY : STD_LOGIC := '0';
SIGNAL BAUD_DIVIDER : INTEGER RANGE 0 TO (FREQUENCY/100 + BAUD/100 - 1) := 0;
BEGIN
	
  	TXD_BUSY <= BUSY; BUSY <= '0' WHEN STATE = IDLE ELSE '1';
	
	BAUD_GEN : PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF BUSY = '1' THEN
				BAUD_DIVIDER <= BAUD_DIVIDER + (BAUD/100);
				IF BAUD_DIVIDER > (FREQUENCY/100) THEN
					BAUD_TICK <= '1';
					BAUD_DIVIDER <= 0;
				ELSE
					BAUD_TICK <= '0';
				END IF;
			END IF;
		END IF;
	END PROCESS BAUD_GEN;

	STATE_PROC : PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			CASE STATE IS
				WHEN IDLE =>
					IF TXD_START = '1' THEN
						STATE <= START;
					END IF;
				WHEN START =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT0;
					END IF;
				WHEN BIT0 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT1;
					END IF;
				WHEN BIT1 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT2;
					END IF;
				WHEN BIT2 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT3;
					END IF;
				WHEN BIT3 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT4;
					END IF;
				WHEN BIT4 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT5;
					END IF;
				WHEN BIT5 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT6;
					END IF;
				WHEN BIT6 =>
					IF BAUD_TICK = '1' THEN
						STATE <= BIT7;
					END IF;
				WHEN BIT7 =>
					IF BAUD_TICK = '1' THEN
						STATE <= STOP1;
					END IF;
				WHEN STOP1 =>
					IF BAUD_TICK = '1' THEN
						STATE <= STOP2;
					END IF;
				WHEN STOP2 =>
					IF BAUD_TICK = '1' THEN
						STATE <= IDLE;
					END IF;
			END CASE;
		END IF;
	END PROCESS STATE_PROC;

	
	DATA_LOAD_PROC : PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF TXD_START = '1' THEN
				DATA <= TXD_DATA;
			END IF;
		END IF;
	END PROCESS DATA_LOAD_PROC;

	
	TXD_PROC : PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			CASE STATE IS
				WHEN IDLE => TXD <= '1';
				WHEN START => TXD <= '0';
				WHEN BIT0 => TXD <= DATA(0);
				WHEN BIT1 => TXD <= DATA(1);
				WHEN BIT2 => TXD <= DATA(2);
				WHEN BIT3 => TXD <= DATA(3);
				WHEN BIT4 => TXD <= DATA(4);
				WHEN BIT5 => TXD <= DATA(5);
				WHEN BIT6 => TXD <= DATA(6);
				WHEN BIT7 => TXD <= DATA(7);
				WHEN STOP1 => TXD <= '1';
				WHEN STOP2 => TXD <= '1';
			END CASE;
		END IF;
	END PROCESS TXD_PROC;

END TRANSMITTER_BEH;


